-- generated with romgen v3.0 by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity bootrom_ab is
	port (
		clk		: in    std_logic;
		addr		: in    std_logic_vector(12 downto 0);
		data		: out   std_logic_vector(7 downto 0)
	);
end;

architecture rtl of bootrom_ab is

	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"F3",x"ED",x"56",x"C3",x"69",x"00",x"00",x"00", -- 0x0000
		x"C3",x"2E",x"00",x"5A",x"38",x"38",x"44",x"4B", -- 0x0008
		x"C3",x"2E",x"00",x"32",x"2E",x"32",x"30",x"00", -- 0x0010
		x"C3",x"2E",x"00",x"1B",x"1B",x"1B",x"C9",x"00", -- 0x0018
		x"C3",x"2E",x"00",x"0B",x"0B",x"0B",x"C9",x"00", -- 0x0020
		x"C3",x"2E",x"00",x"E1",x"E1",x"E1",x"C9",x"00", -- 0x0028
		x"C3",x"2E",x"00",x"FD",x"E9",x"DD",x"E9",x"00", -- 0x0030
		x"C3",x"CD",x"00",x"77",x"23",x"77",x"23",x"77", -- 0x0038
		x"23",x"77",x"23",x"77",x"23",x"77",x"23",x"77", -- 0x0040
		x"23",x"77",x"23",x"77",x"23",x"77",x"23",x"77", -- 0x0048
		x"23",x"77",x"23",x"77",x"23",x"77",x"23",x"77", -- 0x0050
		x"23",x"77",x"23",x"C9",x"23",x"23",x"23",x"23", -- 0x0058
		x"23",x"23",x"23",x"23",x"C9",x"00",x"C3",x"D0", -- 0x0060
		x"00",x"31",x"00",x"00",x"21",x"06",x"14",x"11", -- 0x0068
		x"00",x"5B",x"01",x"06",x"00",x"CD",x"05",x"03", -- 0x0070
		x"21",x"06",x"5B",x"01",x"6E",x"04",x"1E",x"00", -- 0x0078
		x"CD",x"12",x"03",x"CD",x"29",x"0C",x"E5",x"E1", -- 0x0080
		x"76",x"18",x"FE",x"E1",x"E3",x"C3",x"90",x"00", -- 0x0088
		x"7C",x"0F",x"0F",x"0F",x"E6",x"E0",x"B5",x"6F", -- 0x0090
		x"7C",x"E6",x"18",x"F6",x"40",x"67",x"C9",x"7D", -- 0x0098
		x"E6",x"07",x"6F",x"3A",x"00",x"5B",x"E6",x"F8", -- 0x00A0
		x"B5",x"32",x"00",x"5B",x"D3",x"FE",x"C9",x"E1", -- 0x00A8
		x"E1",x"E1",x"E1",x"21",x"00",x"00",x"37",x"C9", -- 0x00B0
		x"E1",x"E1",x"E1",x"2E",x"FF",x"26",x"00",x"22", -- 0x00B8
		x"06",x"5B",x"C3",x"C8",x"00",x"E1",x"E1",x"E1", -- 0x00C0
		x"21",x"FF",x"FF",x"37",x"C9",x"FB",x"ED",x"4D", -- 0x00C8
		x"ED",x"45",x"7B",x"2F",x"5F",x"7A",x"2F",x"57", -- 0x00D0
		x"13",x"C9",x"7D",x"2F",x"6F",x"7C",x"2F",x"67", -- 0x00D8
		x"23",x"C9",x"F1",x"E1",x"D1",x"F5",x"C3",x"FE", -- 0x00E0
		x"00",x"F1",x"E1",x"D1",x"F5",x"CD",x"FE",x"00", -- 0x00E8
		x"EB",x"C9",x"F1",x"D9",x"E1",x"D1",x"D9",x"E1", -- 0x00F0
		x"D1",x"F5",x"C3",x"6A",x"01",x"EB",x"7A",x"B3", -- 0x00F8
		x"28",x"1C",x"44",x"4A",x"C5",x"CB",x"7C",x"C4", -- 0x0100
		x"DA",x"00",x"CB",x"7A",x"C4",x"D2",x"00",x"CD", -- 0x0108
		x"2E",x"01",x"C1",x"78",x"A9",x"FA",x"DA",x"00", -- 0x0110
		x"CB",x"78",x"C8",x"C3",x"D2",x"00",x"EB",x"CD", -- 0x0118
		x"BB",x"00",x"26",x"7F",x"CB",x"7A",x"C8",x"23", -- 0x0120
		x"C9",x"EB",x"7A",x"B3",x"28",x"32",x"14",x"15", -- 0x0128
		x"28",x"1C",x"7D",x"6C",x"26",x"00",x"06",x"08", -- 0x0130
		x"17",x"ED",x"6A",x"ED",x"52",x"30",x"01",x"19", -- 0x0138
		x"3F",x"10",x"F5",x"17",x"50",x"5F",x"EB",x"B7", -- 0x0140
		x"C9",x"EB",x"1C",x"1D",x"28",x"12",x"AF",x"57", -- 0x0148
		x"06",x"10",x"29",x"17",x"38",x"03",x"BB",x"38", -- 0x0150
		x"02",x"93",x"2C",x"10",x"F5",x"5F",x"B7",x"C9", -- 0x0158
		x"EB",x"C3",x"BB",x"00",x"E5",x"D9",x"D1",x"C3", -- 0x0160
		x"D8",x"01",x"AF",x"B3",x"B2",x"D9",x"B3",x"B2", -- 0x0168
		x"28",x"F2",x"E5",x"D9",x"4D",x"44",x"E1",x"D5", -- 0x0170
		x"EB",x"D9",x"C1",x"D5",x"D9",x"C5",x"D5",x"D9", -- 0x0178
		x"C5",x"63",x"69",x"E5",x"D9",x"63",x"69",x"E5", -- 0x0180
		x"62",x"68",x"E5",x"62",x"50",x"69",x"43",x"ED", -- 0x0188
		x"30",x"EB",x"ED",x"30",x"AF",x"19",x"8F",x"59", -- 0x0190
		x"50",x"ED",x"30",x"47",x"4C",x"7A",x"85",x"67", -- 0x0198
		x"6B",x"D1",x"ED",x"30",x"EB",x"ED",x"4A",x"EB", -- 0x01A0
		x"D5",x"D9",x"C1",x"E1",x"D1",x"7C",x"62",x"57", -- 0x01A8
		x"ED",x"30",x"EB",x"ED",x"30",x"09",x"19",x"44", -- 0x01B0
		x"4D",x"E1",x"D1",x"7C",x"62",x"57",x"ED",x"30", -- 0x01B8
		x"EB",x"ED",x"30",x"78",x"83",x"85",x"E1",x"D1", -- 0x01C0
		x"44",x"62",x"50",x"ED",x"30",x"EB",x"ED",x"30", -- 0x01C8
		x"85",x"83",x"47",x"C5",x"D9",x"D1",x"AF",x"C9", -- 0x01D0
		x"45",x"4B",x"5D",x"6A",x"E5",x"69",x"ED",x"30", -- 0x01D8
		x"EB",x"ED",x"30",x"AF",x"19",x"8F",x"59",x"50", -- 0x01E0
		x"ED",x"30",x"47",x"4C",x"7A",x"85",x"67",x"6B", -- 0x01E8
		x"D1",x"ED",x"30",x"EB",x"ED",x"4A",x"EB",x"C9", -- 0x01F0
		x"37",x"C5",x"D9",x"E1",x"11",x"00",x"00",x"D2", -- 0x01F8
		x"0C",x"02",x"C3",x"06",x"02",x"D9",x"7A",x"B3", -- 0x0200
		x"B4",x"B5",x"28",x"42",x"AF",x"E5",x"D9",x"4D", -- 0x0208
		x"44",x"E1",x"D5",x"EB",x"6F",x"67",x"D9",x"C1", -- 0x0210
		x"6F",x"67",x"78",x"06",x"20",x"D9",x"CB",x"11", -- 0x0218
		x"CB",x"10",x"D9",x"CB",x"11",x"17",x"D9",x"ED", -- 0x0220
		x"6A",x"D9",x"ED",x"6A",x"D9",x"ED",x"52",x"D9", -- 0x0228
		x"ED",x"52",x"30",x"05",x"D9",x"19",x"D9",x"ED", -- 0x0230
		x"5A",x"3F",x"10",x"E1",x"D9",x"CB",x"11",x"CB", -- 0x0238
		x"10",x"D9",x"CB",x"11",x"17",x"E5",x"D9",x"D1", -- 0x0240
		x"C5",x"D9",x"E1",x"59",x"57",x"C9",x"1B",x"C3", -- 0x0248
		x"BB",x"00",x"E1",x"D1",x"E3",x"C3",x"58",x"02", -- 0x0250
		x"E5",x"CD",x"D8",x"01",x"01",x"E8",x"03",x"CD", -- 0x0258
		x"F9",x"01",x"C1",x"E5",x"11",x"06",x"00",x"21", -- 0x0260
		x"FC",x"AC",x"CD",x"F9",x"01",x"B7",x"11",x"1E", -- 0x0268
		x"00",x"ED",x"52",x"D1",x"C3",x"77",x"02",x"7A", -- 0x0270
		x"B3",x"C8",x"1B",x"7D",x"CB",x"3D",x"CB",x"3D", -- 0x0278
		x"2F",x"E6",x"03",x"4F",x"06",x"00",x"FD",x"21", -- 0x0280
		x"8F",x"02",x"FD",x"09",x"CD",x"C2",x"02",x"00", -- 0x0288
		x"00",x"00",x"04",x"0C",x"0D",x"20",x"FD",x"0E", -- 0x0290
		x"3F",x"05",x"C2",x"94",x"02",x"EE",x"10",x"D3", -- 0x0298
		x"FE",x"44",x"4F",x"CB",x"67",x"20",x"09",x"7A", -- 0x02A0
		x"B3",x"79",x"28",x"08",x"4D",x"1B",x"FD",x"E9", -- 0x02A8
		x"4D",x"0C",x"FD",x"E9",x"C3",x"B7",x"02",x"4F", -- 0x02B0
		x"3A",x"00",x"5B",x"E6",x"E8",x"B1",x"32",x"00", -- 0x02B8
		x"5B",x"C9",x"3A",x"00",x"5B",x"E6",x"17",x"C9", -- 0x02C0
		x"11",x"0A",x"5B",x"1A",x"B7",x"CA",x"86",x"00", -- 0x02C8
		x"E5",x"6F",x"26",x"00",x"29",x"19",x"47",x"56", -- 0x02D0
		x"2B",x"5E",x"2B",x"C5",x"E5",x"EB",x"CD",x"34", -- 0x02D8
		x"00",x"E1",x"C1",x"10",x"F2",x"E1",x"C3",x"86", -- 0x02E0
		x"00",x"F1",x"D1",x"E1",x"C1",x"F5",x"C3",x"F1", -- 0x02E8
		x"02",x"78",x"B1",x"28",x"09",x"1A",x"ED",x"A1", -- 0x02F0
		x"20",x"07",x"13",x"EA",x"F5",x"02",x"60",x"69", -- 0x02F8
		x"C9",x"2B",x"96",x"67",x"C9",x"78",x"B1",x"28", -- 0x0300
		x"06",x"D5",x"ED",x"B0",x"E1",x"B7",x"C9",x"62", -- 0x0308
		x"6B",x"C9",x"78",x"B1",x"7B",x"54",x"5D",x"C8", -- 0x0310
		x"77",x"13",x"0B",x"78",x"B1",x"C8",x"E5",x"ED", -- 0x0318
		x"B0",x"E1",x"C9",x"AF",x"4F",x"47",x"ED",x"B1", -- 0x0320
		x"21",x"FF",x"FF",x"ED",x"42",x"C9",x"5D",x"54", -- 0x0328
		x"1B",x"7A",x"B3",x"28",x"08",x"21",x"81",x"0D", -- 0x0330
		x"CD",x"43",x"03",x"18",x"F3",x"21",x"76",x"0D", -- 0x0338
		x"C3",x"43",x"03",x"01",x"73",x"FF",x"09",x"01", -- 0x0340
		x"E9",x"FF",x"09",x"38",x"FD",x"7D",x"C6",x"0F", -- 0x0348
		x"30",x"06",x"FE",x"08",x"38",x"03",x"F6",x"00", -- 0x0350
		x"23",x"1F",x"38",x"01",x"00",x"1F",x"30",x"02", -- 0x0358
		x"F6",x"00",x"1F",x"D0",x"C9",x"DD",x"E5",x"DD", -- 0x0360
		x"21",x"00",x"00",x"DD",x"39",x"3A",x"0C",x"5B", -- 0x0368
		x"B7",x"28",x"36",x"DD",x"6E",x"04",x"DD",x"66", -- 0x0370
		x"05",x"22",x"3C",x"5D",x"DD",x"6E",x"06",x"DD", -- 0x0378
		x"66",x"07",x"22",x"3E",x"5D",x"06",x"07",x"21", -- 0x0380
		x"3F",x"5D",x"CB",x"3E",x"2B",x"CB",x"1E",x"2B", -- 0x0388
		x"CB",x"1E",x"2B",x"CB",x"1E",x"10",x"F0",x"DD", -- 0x0390
		x"7E",x"04",x"E6",x"7F",x"21",x"38",x"5D",x"77", -- 0x0398
		x"AF",x"23",x"77",x"23",x"77",x"23",x"77",x"18", -- 0x03A0
		x"22",x"DD",x"6E",x"05",x"DD",x"66",x"06",x"22", -- 0x03A8
		x"3C",x"5D",x"21",x"3D",x"5D",x"DD",x"7E",x"07", -- 0x03B0
		x"23",x"77",x"23",x"36",x"00",x"DD",x"7E",x"04", -- 0x03B8
		x"21",x"38",x"5D",x"77",x"AF",x"23",x"77",x"23", -- 0x03C0
		x"77",x"23",x"77",x"2A",x"3C",x"5D",x"ED",x"4B", -- 0x03C8
		x"34",x"5D",x"AF",x"ED",x"42",x"20",x"10",x"3A", -- 0x03D0
		x"3E",x"5D",x"21",x"36",x"5D",x"96",x"20",x"07", -- 0x03D8
		x"3A",x"3F",x"5D",x"23",x"96",x"28",x"43",x"2A", -- 0x03E0
		x"0D",x"5B",x"ED",x"4B",x"3C",x"5D",x"09",x"3A", -- 0x03E8
		x"0F",x"5B",x"4D",x"44",x"21",x"3E",x"5D",x"8E", -- 0x03F0
		x"5F",x"3A",x"10",x"5B",x"21",x"3F",x"5D",x"8E", -- 0x03F8
		x"57",x"21",x"33",x"5B",x"E5",x"D5",x"C5",x"CD", -- 0x0400
		x"6B",x"0F",x"7D",x"B7",x"20",x"07",x"21",x"00", -- 0x0408
		x"00",x"5D",x"55",x"18",x"4F",x"21",x"3C",x"5D", -- 0x0410
		x"7E",x"EB",x"21",x"34",x"5D",x"77",x"23",x"13", -- 0x0418
		x"1A",x"77",x"23",x"13",x"1A",x"77",x"23",x"13", -- 0x0420
		x"1A",x"77",x"ED",x"4B",x"38",x"5D",x"3A",x"0C", -- 0x0428
		x"5B",x"B7",x"28",x"15",x"69",x"60",x"29",x"29", -- 0x0430
		x"11",x"33",x"5B",x"19",x"4E",x"23",x"46",x"23", -- 0x0438
		x"5E",x"23",x"7E",x"6B",x"E6",x"0F",x"67",x"18", -- 0x0440
		x"0D",x"11",x"33",x"5B",x"69",x"60",x"29",x"19", -- 0x0448
		x"4E",x"23",x"46",x"21",x"00",x"00",x"ED",x"43", -- 0x0450
		x"38",x"5D",x"22",x"3A",x"5D",x"2A",x"38",x"5D", -- 0x0458
		x"ED",x"5B",x"3A",x"5D",x"DD",x"E1",x"C9",x"DD", -- 0x0460
		x"E5",x"DD",x"21",x"00",x"00",x"DD",x"39",x"21", -- 0x0468
		x"F8",x"FF",x"39",x"F9",x"21",x"FF",x"FF",x"22", -- 0x0470
		x"34",x"5D",x"22",x"36",x"5D",x"21",x"0C",x"5B", -- 0x0478
		x"36",x"00",x"21",x"33",x"5B",x"E5",x"21",x"00", -- 0x0480
		x"00",x"E5",x"E5",x"CD",x"6B",x"0F",x"7D",x"B7", -- 0x0488
		x"20",x"04",x"6F",x"C3",x"77",x"08",x"21",x"00", -- 0x0490
		x"00",x"22",x"40",x"5D",x"22",x"42",x"5D",x"21", -- 0x0498
		x"33",x"5D",x"36",x"01",x"21",x"08",x"00",x"E5", -- 0x04A0
		x"21",x"2B",x"13",x"E5",x"21",x"69",x"5B",x"E5", -- 0x04A8
		x"CD",x"E9",x"02",x"7C",x"B5",x"20",x"05",x"21", -- 0x04B0
		x"33",x"5D",x"36",x"00",x"21",x"08",x"00",x"E5", -- 0x04B8
		x"21",x"34",x"13",x"E5",x"21",x"85",x"5B",x"E5", -- 0x04C0
		x"CD",x"E9",x"02",x"7C",x"B5",x"20",x"05",x"21", -- 0x04C8
		x"33",x"5D",x"36",x"00",x"3A",x"33",x"5D",x"B7", -- 0x04D0
		x"28",x"63",x"21",x"33",x"5B",x"22",x"44",x"5D", -- 0x04D8
		x"ED",x"4B",x"44",x"5D",x"21",x"C6",x"01",x"09", -- 0x04E0
		x"E5",x"11",x"40",x"5D",x"ED",x"A0",x"03",x"ED", -- 0x04E8
		x"A0",x"03",x"ED",x"A0",x"03",x"7E",x"12",x"D1", -- 0x04F0
		x"21",x"FE",x"01",x"09",x"7E",x"23",x"46",x"4F", -- 0x04F8
		x"D6",x"AA",x"20",x"13",x"78",x"D6",x"55",x"20", -- 0x0500
		x"0E",x"EB",x"11",x"40",x"5D",x"ED",x"A0",x"ED", -- 0x0508
		x"A0",x"ED",x"A0",x"7E",x"12",x"18",x"0F",x"79", -- 0x0510
		x"D6",x"55",x"20",x"05",x"78",x"D6",x"AA",x"28", -- 0x0518
		x"05",x"2E",x"00",x"C3",x"77",x"08",x"21",x"33", -- 0x0520
		x"5B",x"E5",x"2A",x"42",x"5D",x"E5",x"2A",x"40", -- 0x0528
		x"5D",x"E5",x"CD",x"6B",x"0F",x"7D",x"B7",x"20", -- 0x0530
		x"04",x"6F",x"C3",x"77",x"08",x"21",x"08",x"00", -- 0x0538
		x"E5",x"21",x"34",x"13",x"E5",x"21",x"85",x"5B", -- 0x0540
		x"E5",x"CD",x"E9",x"02",x"7C",x"B5",x"20",x"07", -- 0x0548
		x"21",x"0C",x"5B",x"36",x"01",x"18",x"18",x"21", -- 0x0550
		x"08",x"00",x"E5",x"21",x"2B",x"13",x"E5",x"21", -- 0x0558
		x"69",x"5B",x"E5",x"CD",x"E9",x"02",x"7C",x"B5", -- 0x0560
		x"28",x"05",x"2E",x"00",x"C3",x"77",x"08",x"3A", -- 0x0568
		x"31",x"5D",x"D6",x"55",x"20",x"07",x"3A",x"32", -- 0x0570
		x"5D",x"D6",x"AA",x"28",x"05",x"2E",x"00",x"C3", -- 0x0578
		x"77",x"08",x"3A",x"33",x"5B",x"FE",x"E9",x"28", -- 0x0580
		x"09",x"D6",x"EB",x"28",x"05",x"2E",x"00",x"C3", -- 0x0588
		x"77",x"08",x"3A",x"3E",x"5B",x"B7",x"20",x"07", -- 0x0590
		x"3A",x"3F",x"5B",x"D6",x"02",x"28",x"05",x"2E", -- 0x0598
		x"00",x"C3",x"77",x"08",x"3A",x"40",x"5B",x"21", -- 0x05A0
		x"23",x"5B",x"77",x"AF",x"23",x"77",x"23",x"77", -- 0x05A8
		x"23",x"77",x"2A",x"23",x"5B",x"01",x"FF",x"FF", -- 0x05B0
		x"09",x"22",x"27",x"5B",x"3A",x"25",x"5B",x"CE", -- 0x05B8
		x"FF",x"32",x"29",x"5B",x"3A",x"26",x"5B",x"CE", -- 0x05C0
		x"FF",x"32",x"2A",x"5B",x"3A",x"41",x"5B",x"4F", -- 0x05C8
		x"11",x"00",x"00",x"43",x"21",x"40",x"5D",x"7E", -- 0x05D0
		x"81",x"DD",x"77",x"FC",x"23",x"7E",x"88",x"DD", -- 0x05D8
		x"77",x"FD",x"23",x"7E",x"8B",x"DD",x"77",x"FE", -- 0x05E0
		x"23",x"7E",x"8A",x"DD",x"77",x"FF",x"3A",x"42", -- 0x05E8
		x"5B",x"0E",x"00",x"47",x"11",x"00",x"00",x"DD", -- 0x05F0
		x"7E",x"FC",x"81",x"21",x"0D",x"5B",x"77",x"DD", -- 0x05F8
		x"7E",x"FD",x"88",x"23",x"77",x"DD",x"7E",x"FE", -- 0x0600
		x"8B",x"23",x"77",x"DD",x"7E",x"FF",x"8A",x"23", -- 0x0608
		x"77",x"3A",x"43",x"5B",x"6F",x"26",x"00",x"22", -- 0x0610
		x"21",x"5B",x"3A",x"0C",x"5B",x"B7",x"CA",x"C2", -- 0x0618
		x"07",x"21",x"08",x"00",x"E5",x"21",x"34",x"13", -- 0x0620
		x"E5",x"21",x"85",x"5B",x"E5",x"CD",x"E9",x"02", -- 0x0628
		x"7C",x"B5",x"28",x"05",x"2E",x"00",x"C3",x"77", -- 0x0630
		x"08",x"2A",x"23",x"5B",x"22",x"2B",x"5B",x"2A", -- 0x0638
		x"25",x"5B",x"22",x"2D",x"5B",x"06",x"04",x"21", -- 0x0640
		x"2B",x"5B",x"CB",x"26",x"23",x"CB",x"16",x"23", -- 0x0648
		x"CB",x"16",x"23",x"CB",x"16",x"10",x"F0",x"21", -- 0x0650
		x"23",x"5B",x"7E",x"EB",x"21",x"1D",x"5B",x"77", -- 0x0658
		x"23",x"13",x"1A",x"77",x"23",x"13",x"1A",x"77", -- 0x0660
		x"23",x"13",x"1A",x"77",x"3A",x"57",x"5B",x"21", -- 0x0668
		x"58",x"5B",x"4E",x"11",x"00",x"00",x"DD",x"71", -- 0x0670
		x"FD",x"DD",x"73",x"FE",x"DD",x"73",x"FF",x"DD", -- 0x0678
		x"36",x"FC",x"00",x"01",x"00",x"00",x"1E",x"00", -- 0x0680
		x"DD",x"86",x"FC",x"DD",x"77",x"F8",x"79",x"DD", -- 0x0688
		x"8E",x"FD",x"DD",x"77",x"F9",x"78",x"DD",x"8E", -- 0x0690
		x"FE",x"DD",x"77",x"FA",x"7B",x"DD",x"8E",x"FF", -- 0x0698
		x"DD",x"77",x"FB",x"3A",x"59",x"5B",x"0E",x"00", -- 0x06A0
		x"57",x"AF",x"5F",x"DD",x"86",x"F8",x"DD",x"77", -- 0x06A8
		x"FC",x"7B",x"DD",x"8E",x"F9",x"DD",x"77",x"FD", -- 0x06B0
		x"7A",x"DD",x"8E",x"FA",x"DD",x"77",x"FE",x"79", -- 0x06B8
		x"DD",x"8E",x"FB",x"DD",x"77",x"FF",x"3A",x"5A", -- 0x06C0
		x"5B",x"4F",x"11",x"00",x"00",x"43",x"DD",x"7E", -- 0x06C8
		x"FC",x"80",x"21",x"2F",x"5B",x"77",x"DD",x"7E", -- 0x06D0
		x"FD",x"8B",x"23",x"77",x"DD",x"7E",x"FE",x"8A", -- 0x06D8
		x"23",x"77",x"DD",x"7E",x"FF",x"89",x"23",x"77", -- 0x06E0
		x"ED",x"4B",x"21",x"5B",x"11",x"00",x"00",x"2A", -- 0x06E8
		x"31",x"5B",x"E5",x"2A",x"2F",x"5B",x"E5",x"D5", -- 0x06F0
		x"C5",x"CD",x"F2",x"00",x"ED",x"4B",x"0D",x"5B", -- 0x06F8
		x"09",x"22",x"11",x"5B",x"2A",x"0F",x"5B",x"ED", -- 0x0700
		x"5A",x"22",x"13",x"5B",x"3A",x"5F",x"5B",x"21", -- 0x0708
		x"60",x"5B",x"4E",x"11",x"00",x"00",x"DD",x"71", -- 0x0710
		x"FD",x"DD",x"73",x"FE",x"DD",x"73",x"FF",x"DD", -- 0x0718
		x"36",x"FC",x"00",x"01",x"00",x"00",x"1E",x"00", -- 0x0720
		x"DD",x"86",x"FC",x"DD",x"77",x"F8",x"79",x"DD", -- 0x0728
		x"8E",x"FD",x"DD",x"77",x"F9",x"78",x"DD",x"8E", -- 0x0730
		x"FE",x"DD",x"77",x"FA",x"7B",x"DD",x"8E",x"FF", -- 0x0738
		x"DD",x"77",x"FB",x"3A",x"61",x"5B",x"0E",x"00", -- 0x0740
		x"57",x"AF",x"5F",x"DD",x"86",x"F8",x"DD",x"77", -- 0x0748
		x"FC",x"7B",x"DD",x"8E",x"F9",x"DD",x"77",x"FD", -- 0x0750
		x"7A",x"DD",x"8E",x"FA",x"DD",x"77",x"FE",x"79", -- 0x0758
		x"DD",x"8E",x"FB",x"DD",x"77",x"FF",x"3A",x"62", -- 0x0760
		x"5B",x"E6",x"0F",x"0E",x"00",x"47",x"79",x"07", -- 0x0768
		x"ED",x"62",x"11",x"00",x"00",x"4B",x"DD",x"7E", -- 0x0770
		x"FC",x"81",x"21",x"15",x"5B",x"77",x"DD",x"7E", -- 0x0778
		x"FD",x"8B",x"23",x"77",x"DD",x"7E",x"FE",x"8A", -- 0x0780
		x"23",x"77",x"DD",x"7E",x"FF",x"88",x"23",x"77", -- 0x0788
		x"2A",x"15",x"5B",x"01",x"FE",x"FF",x"09",x"4D", -- 0x0790
		x"44",x"2A",x"17",x"5B",x"11",x"FF",x"FF",x"ED", -- 0x0798
		x"5A",x"EB",x"2A",x"25",x"5B",x"E5",x"2A",x"23", -- 0x07A0
		x"5B",x"E5",x"D5",x"C5",x"CD",x"F2",x"00",x"ED", -- 0x07A8
		x"4B",x"11",x"5B",x"09",x"22",x"19",x"5B",x"2A", -- 0x07B0
		x"13",x"5B",x"ED",x"5A",x"22",x"1B",x"5B",x"C3", -- 0x07B8
		x"75",x"08",x"3A",x"44",x"5B",x"06",x"00",x"21", -- 0x07C0
		x"45",x"5B",x"66",x"2E",x"00",x"4F",x"09",x"22", -- 0x07C8
		x"2B",x"5B",x"21",x"00",x"00",x"22",x"2D",x"5B", -- 0x07D0
		x"21",x"2B",x"5B",x"7E",x"23",x"4E",x"23",x"5E", -- 0x07D8
		x"23",x"56",x"06",x"05",x"87",x"CB",x"11",x"CB", -- 0x07E0
		x"13",x"CB",x"12",x"10",x"F7",x"C6",x"FF",x"79", -- 0x07E8
		x"CE",x"01",x"4F",x"30",x"01",x"13",x"21",x"1D", -- 0x07F0
		x"5B",x"71",x"23",x"73",x"23",x"72",x"23",x"36", -- 0x07F8
		x"00",x"2B",x"CB",x"3E",x"2B",x"CB",x"1E",x"2B", -- 0x0800
		x"CB",x"1E",x"3A",x"49",x"5B",x"06",x"00",x"21", -- 0x0808
		x"4A",x"5B",x"66",x"2E",x"00",x"4F",x"09",x"22", -- 0x0810
		x"2F",x"5B",x"21",x"00",x"00",x"22",x"31",x"5B", -- 0x0818
		x"ED",x"4B",x"21",x"5B",x"11",x"00",x"00",x"2A", -- 0x0820
		x"31",x"5B",x"E5",x"2A",x"2F",x"5B",x"E5",x"D5", -- 0x0828
		x"C5",x"CD",x"F2",x"00",x"ED",x"4B",x"0D",x"5B", -- 0x0830
		x"09",x"22",x"19",x"5B",x"2A",x"0F",x"5B",x"ED", -- 0x0838
		x"5A",x"22",x"1B",x"5B",x"21",x"00",x"00",x"22", -- 0x0840
		x"15",x"5B",x"22",x"17",x"5B",x"3A",x"19",x"5B", -- 0x0848
		x"21",x"1D",x"5B",x"86",x"32",x"11",x"5B",x"3A", -- 0x0850
		x"1A",x"5B",x"21",x"1E",x"5B",x"8E",x"32",x"12", -- 0x0858
		x"5B",x"3A",x"1B",x"5B",x"21",x"1F",x"5B",x"8E", -- 0x0860
		x"32",x"13",x"5B",x"3A",x"1C",x"5B",x"21",x"20", -- 0x0868
		x"5B",x"8E",x"32",x"14",x"5B",x"2E",x"01",x"DD", -- 0x0870
		x"F9",x"DD",x"E1",x"C9",x"DD",x"E5",x"DD",x"21", -- 0x0878
		x"00",x"00",x"DD",x"39",x"21",x"F8",x"FF",x"39", -- 0x0880
		x"F9",x"21",x"00",x"00",x"22",x"46",x"5D",x"22", -- 0x0888
		x"48",x"5D",x"AF",x"6F",x"67",x"22",x"4A",x"5D", -- 0x0890
		x"21",x"FF",x"FF",x"22",x"34",x"5D",x"22",x"36", -- 0x0898
		x"5D",x"21",x"15",x"5B",x"7E",x"EB",x"21",x"50", -- 0x08A0
		x"5D",x"77",x"23",x"13",x"1A",x"77",x"23",x"13", -- 0x08A8
		x"1A",x"77",x"23",x"13",x"1A",x"77",x"21",x"19", -- 0x08B0
		x"5B",x"7E",x"EB",x"21",x"4C",x"5D",x"77",x"23", -- 0x08B8
		x"13",x"1A",x"77",x"23",x"13",x"1A",x"77",x"23", -- 0x08C0
		x"13",x"1A",x"77",x"3A",x"0C",x"5B",x"B7",x"28", -- 0x08C8
		x"17",x"21",x"23",x"5B",x"7E",x"23",x"4E",x"23", -- 0x08D0
		x"5E",x"23",x"56",x"06",x"04",x"87",x"CB",x"11", -- 0x08D8
		x"CB",x"13",x"CB",x"12",x"10",x"F7",x"18",x"15", -- 0x08E0
		x"21",x"1D",x"5B",x"7E",x"23",x"4E",x"23",x"5E", -- 0x08E8
		x"23",x"56",x"06",x"04",x"87",x"CB",x"11",x"CB", -- 0x08F0
		x"13",x"CB",x"12",x"10",x"F7",x"21",x"58",x"5D", -- 0x08F8
		x"77",x"23",x"71",x"23",x"73",x"23",x"72",x"21", -- 0x0900
		x"00",x"00",x"22",x"54",x"5D",x"22",x"56",x"5D", -- 0x0908
		x"2A",x"54",x"5D",x"ED",x"4B",x"58",x"5D",x"AF", -- 0x0910
		x"ED",x"42",x"20",x"11",x"3A",x"56",x"5D",x"21", -- 0x0918
		x"5A",x"5D",x"96",x"20",x"08",x"3A",x"57",x"5D", -- 0x0920
		x"23",x"96",x"CA",x"57",x"0A",x"3A",x"54",x"5D", -- 0x0928
		x"E6",x"0F",x"20",x"29",x"ED",x"4B",x"4C",x"5D", -- 0x0930
		x"ED",x"5B",x"4E",x"5D",x"21",x"4C",x"5D",x"34", -- 0x0938
		x"20",x"0A",x"23",x"34",x"20",x"06",x"23",x"34", -- 0x0940
		x"20",x"02",x"23",x"34",x"21",x"33",x"5B",x"E5", -- 0x0948
		x"D5",x"C5",x"CD",x"6B",x"0F",x"21",x"33",x"5B", -- 0x0950
		x"22",x"4A",x"5D",x"18",x"0A",x"2A",x"4A",x"5D", -- 0x0958
		x"11",x"20",x"00",x"19",x"22",x"4A",x"5D",x"ED", -- 0x0960
		x"4B",x"4A",x"5D",x"0A",x"B7",x"CA",x"41",x"0A", -- 0x0968
		x"D6",x"E5",x"CA",x"41",x"0A",x"21",x"0B",x"00", -- 0x0970
		x"09",x"7E",x"E6",x"18",x"C2",x"41",x"0A",x"DD", -- 0x0978
		x"5E",x"06",x"DD",x"56",x"07",x"21",x"0B",x"00", -- 0x0980
		x"E5",x"D5",x"C5",x"CD",x"E9",x"02",x"7C",x"B5", -- 0x0988
		x"C2",x"41",x"0A",x"DD",x"7E",x"04",x"DD",x"77", -- 0x0990
		x"F8",x"DD",x"7E",x"05",x"DD",x"77",x"F9",x"DD", -- 0x0998
		x"7E",x"F8",x"C6",x"04",x"5F",x"DD",x"7E",x"F9", -- 0x09A0
		x"CE",x"00",x"57",x"2A",x"4A",x"5D",x"D5",x"EB", -- 0x09A8
		x"21",x"06",x"00",x"39",x"EB",x"01",x"1C",x"00", -- 0x09B0
		x"09",x"01",x"04",x"00",x"ED",x"B0",x"D1",x"21", -- 0x09B8
		x"04",x"00",x"39",x"01",x"04",x"00",x"ED",x"B0", -- 0x09C0
		x"DD",x"7E",x"F8",x"C6",x"08",x"DD",x"77",x"FA", -- 0x09C8
		x"DD",x"7E",x"F9",x"CE",x"00",x"DD",x"77",x"FB", -- 0x09D0
		x"ED",x"4B",x"4A",x"5D",x"21",x"1A",x"00",x"09", -- 0x09D8
		x"5E",x"23",x"56",x"3A",x"0C",x"5B",x"B7",x"28", -- 0x09E0
		x"18",x"21",x"14",x"00",x"09",x"46",x"23",x"7E", -- 0x09E8
		x"E6",x"0F",x"DD",x"70",x"FE",x"DD",x"77",x"FF", -- 0x09F0
		x"AF",x"DD",x"77",x"FC",x"DD",x"77",x"FD",x"18", -- 0x09F8
		x"0D",x"AF",x"DD",x"77",x"FC",x"DD",x"77",x"FD", -- 0x0A00
		x"DD",x"77",x"FE",x"DD",x"77",x"FF",x"7B",x"01", -- 0x0A08
		x"00",x"00",x"DD",x"86",x"FC",x"5F",x"7A",x"DD", -- 0x0A10
		x"8E",x"FD",x"57",x"79",x"DD",x"8E",x"FE",x"4F", -- 0x0A18
		x"78",x"DD",x"8E",x"FF",x"47",x"DD",x"6E",x"FA", -- 0x0A20
		x"DD",x"66",x"FB",x"73",x"23",x"72",x"23",x"71", -- 0x0A28
		x"23",x"70",x"E1",x"E5",x"AF",x"77",x"23",x"77", -- 0x0A30
		x"23",x"77",x"23",x"77",x"2E",x"01",x"C3",x"C2", -- 0x0A38
		x"0A",x"21",x"54",x"5D",x"34",x"C2",x"10",x"09", -- 0x0A40
		x"23",x"34",x"C2",x"10",x"09",x"23",x"34",x"C2", -- 0x0A48
		x"10",x"09",x"23",x"34",x"C3",x"10",x"09",x"3A", -- 0x0A50
		x"0C",x"5B",x"B7",x"28",x"63",x"2A",x"52",x"5D", -- 0x0A58
		x"E5",x"2A",x"50",x"5D",x"E5",x"CD",x"65",x"03", -- 0x0A60
		x"F1",x"F1",x"22",x"50",x"5D",x"EB",x"22",x"52", -- 0x0A68
		x"5D",x"3A",x"50",x"5D",x"E6",x"F8",x"4F",x"2A", -- 0x0A70
		x"51",x"5D",x"3A",x"53",x"5D",x"E6",x"0F",x"47", -- 0x0A78
		x"79",x"D6",x"F8",x"20",x"0A",x"7D",x"A4",x"3C", -- 0x0A80
		x"20",x"05",x"78",x"D6",x"0F",x"28",x"31",x"2A", -- 0x0A88
		x"50",x"5D",x"01",x"FE",x"FF",x"09",x"4D",x"44", -- 0x0A90
		x"2A",x"52",x"5D",x"11",x"FF",x"FF",x"ED",x"5A", -- 0x0A98
		x"E5",x"C5",x"2A",x"25",x"5B",x"E5",x"2A",x"23", -- 0x0AA0
		x"5B",x"E5",x"CD",x"F2",x"00",x"ED",x"4B",x"11", -- 0x0AA8
		x"5B",x"09",x"22",x"4C",x"5D",x"2A",x"13",x"5B", -- 0x0AB0
		x"ED",x"5A",x"22",x"4E",x"5D",x"C3",x"07",x"09", -- 0x0AB8
		x"2E",x"00",x"DD",x"F9",x"DD",x"E1",x"C9",x"DD", -- 0x0AC0
		x"E5",x"DD",x"21",x"00",x"00",x"DD",x"39",x"F5", -- 0x0AC8
		x"F5",x"21",x"11",x"5B",x"7E",x"EB",x"21",x"5C", -- 0x0AD0
		x"5D",x"77",x"23",x"13",x"1A",x"77",x"23",x"13", -- 0x0AD8
		x"1A",x"77",x"23",x"13",x"1A",x"77",x"DD",x"7E", -- 0x0AE0
		x"04",x"DD",x"77",x"FC",x"6F",x"DD",x"7E",x"05", -- 0x0AE8
		x"DD",x"77",x"FD",x"67",x"11",x"08",x"00",x"19", -- 0x0AF0
		x"DD",x"75",x"FE",x"DD",x"74",x"FF",x"4E",x"23", -- 0x0AF8
		x"46",x"23",x"5E",x"23",x"56",x"21",x"FE",x"FF", -- 0x0B00
		x"09",x"4D",x"44",x"21",x"FF",x"FF",x"ED",x"5A", -- 0x0B08
		x"E5",x"C5",x"2A",x"25",x"5B",x"E5",x"2A",x"23", -- 0x0B10
		x"5B",x"E5",x"CD",x"F2",x"00",x"ED",x"4B",x"5C", -- 0x0B18
		x"5D",x"09",x"22",x"5C",x"5D",x"2A",x"5E",x"5D", -- 0x0B20
		x"ED",x"5A",x"22",x"5E",x"5D",x"E1",x"4E",x"E5", -- 0x0B28
		x"23",x"46",x"23",x"5E",x"23",x"56",x"2A",x"27", -- 0x0B30
		x"5B",x"79",x"A5",x"4F",x"78",x"A4",x"47",x"2A", -- 0x0B38
		x"29",x"5B",x"7B",x"A5",x"5F",x"7A",x"A4",x"57", -- 0x0B40
		x"2A",x"5C",x"5D",x"09",x"22",x"5C",x"5D",x"2A", -- 0x0B48
		x"5E",x"5D",x"ED",x"5A",x"22",x"5E",x"5D",x"DD", -- 0x0B50
		x"6E",x"06",x"DD",x"66",x"07",x"E5",x"2A",x"5E", -- 0x0B58
		x"5D",x"E5",x"2A",x"5C",x"5D",x"E5",x"CD",x"6B", -- 0x0B60
		x"0F",x"7D",x"B7",x"20",x"03",x"6F",x"18",x"54", -- 0x0B68
		x"E1",x"4E",x"E5",x"23",x"46",x"23",x"5E",x"23", -- 0x0B70
		x"56",x"0C",x"20",x"04",x"04",x"20",x"01",x"13", -- 0x0B78
		x"E1",x"E5",x"71",x"23",x"70",x"23",x"73",x"23", -- 0x0B80
		x"72",x"79",x"21",x"27",x"5B",x"A6",x"4F",x"78", -- 0x0B88
		x"23",x"A6",x"47",x"7B",x"23",x"A6",x"5F",x"7A", -- 0x0B90
		x"23",x"A6",x"B3",x"B0",x"B1",x"20",x"23",x"DD", -- 0x0B98
		x"6E",x"FE",x"DD",x"66",x"FF",x"4E",x"23",x"46", -- 0x0BA0
		x"23",x"5E",x"23",x"56",x"D5",x"C5",x"CD",x"65", -- 0x0BA8
		x"03",x"F1",x"F1",x"4D",x"DD",x"6E",x"FE",x"44", -- 0x0BB0
		x"DD",x"66",x"FF",x"71",x"23",x"70",x"23",x"73", -- 0x0BB8
		x"23",x"72",x"2E",x"01",x"DD",x"F9",x"DD",x"E1", -- 0x0BC0
		x"C9",x"DD",x"E5",x"DD",x"21",x"00",x"00",x"DD", -- 0x0BC8
		x"39",x"3E",x"FF",x"D3",x"E7",x"2E",x"02",x"CD", -- 0x0BD0
		x"9F",x"00",x"DD",x"6E",x"04",x"DD",x"66",x"05", -- 0x0BD8
		x"CD",x"23",x"03",x"CB",x"3C",x"CB",x"1D",x"3E", -- 0x0BE0
		x"10",x"95",x"26",x"0C",x"6F",x"E5",x"CD",x"62", -- 0x0BE8
		x"0E",x"F1",x"DD",x"6E",x"04",x"DD",x"66",x"05", -- 0x0BF0
		x"E5",x"CD",x"C2",x"0E",x"F1",x"21",x"FA",x"00", -- 0x0BF8
		x"CD",x"2E",x"03",x"0E",x"00",x"DD",x"7E",x"06", -- 0x0C00
		x"91",x"28",x"15",x"C5",x"21",x"FA",x"00",x"CD", -- 0x0C08
		x"2E",x"03",x"21",x"6E",x"00",x"E5",x"2E",x"7D", -- 0x0C10
		x"E5",x"CD",x"52",x"02",x"C1",x"0C",x"18",x"E5", -- 0x0C18
		x"21",x"01",x"00",x"CD",x"C8",x"02",x"DD",x"E1", -- 0x0C20
		x"C9",x"2E",x"00",x"CD",x"9F",x"00",x"21",x"00", -- 0x0C28
		x"40",x"36",x"00",x"5D",x"54",x"13",x"01",x"FF", -- 0x0C30
		x"17",x"ED",x"B0",x"21",x"00",x"58",x"36",x"07", -- 0x0C38
		x"5D",x"54",x"13",x"01",x"FF",x"02",x"ED",x"B0", -- 0x0C40
		x"CD",x"31",x"0E",x"21",x"B8",x"01",x"E5",x"2E", -- 0x0C48
		x"2C",x"E5",x"CD",x"52",x"02",x"21",x"6C",x"5F", -- 0x0C50
		x"36",x"FA",x"3A",x"6C",x"5F",x"B7",x"28",x"5B", -- 0x0C58
		x"2E",x"10",x"01",x"3B",x"24",x"ED",x"69",x"04", -- 0x0C60
		x"ED",x"68",x"7D",x"E6",x"03",x"3D",x"B7",x"20", -- 0x0C68
		x"4A",x"11",x"0F",x"0C",x"D5",x"CD",x"62",x"0E", -- 0x0C70
		x"F1",x"3A",x"6C",x"5F",x"4F",x"06",x"00",x"21", -- 0x0C78
		x"64",x"00",x"E5",x"C5",x"CD",x"E2",x"00",x"7D", -- 0x0C80
		x"C6",x"30",x"F5",x"33",x"CD",x"83",x"0E",x"33", -- 0x0C88
		x"3A",x"6C",x"5F",x"4F",x"06",x"00",x"21",x"0A", -- 0x0C90
		x"00",x"E5",x"C5",x"CD",x"E2",x"00",x"11",x"0A", -- 0x0C98
		x"00",x"D5",x"E5",x"CD",x"E9",x"00",x"7D",x"C6", -- 0x0CA0
		x"30",x"F5",x"33",x"CD",x"83",x"0E",x"33",x"21", -- 0x0CA8
		x"64",x"00",x"CD",x"2E",x"03",x"21",x"6C",x"5F", -- 0x0CB0
		x"35",x"18",x"9F",x"21",x"00",x"40",x"36",x"00", -- 0x0CB8
		x"5D",x"54",x"13",x"01",x"FF",x"17",x"ED",x"B0", -- 0x0CC0
		x"21",x"00",x"58",x"36",x"02",x"5D",x"54",x"13", -- 0x0CC8
		x"01",x"FF",x"02",x"ED",x"B0",x"21",x"6C",x"5F", -- 0x0CD0
		x"36",x"03",x"CD",x"E2",x"0E",x"7D",x"B7",x"28", -- 0x0CD8
		x"07",x"CD",x"67",x"04",x"7D",x"B7",x"20",x"0C", -- 0x0CE0
		x"21",x"0A",x"00",x"CD",x"2E",x"03",x"21",x"6C", -- 0x0CE8
		x"5F",x"35",x"20",x"E6",x"3A",x"6C",x"5F",x"B7", -- 0x0CF0
		x"20",x"0D",x"3E",x"01",x"F5",x"33",x"21",x"3D", -- 0x0CF8
		x"13",x"E5",x"CD",x"C9",x"0B",x"F1",x"33",x"21", -- 0x0D00
		x"54",x"13",x"E5",x"21",x"60",x"5D",x"E5",x"CD", -- 0x0D08
		x"7C",x"08",x"F1",x"F1",x"7D",x"B7",x"20",x"0D", -- 0x0D10
		x"3E",x"02",x"F5",x"33",x"21",x"60",x"13",x"E5", -- 0x0D18
		x"CD",x"C9",x"0B",x"F1",x"33",x"2E",x"10",x"01", -- 0x0D20
		x"3B",x"24",x"ED",x"69",x"04",x"ED",x"68",x"7D", -- 0x0D28
		x"E6",x"03",x"06",x"00",x"D6",x"03",x"B0",x"C2", -- 0x0D30
		x"15",x"0E",x"21",x"74",x"13",x"E5",x"21",x"60", -- 0x0D38
		x"5D",x"E5",x"CD",x"7C",x"08",x"F1",x"F1",x"7D", -- 0x0D40
		x"B7",x"20",x"0D",x"3E",x"03",x"F5",x"33",x"21", -- 0x0D48
		x"80",x"13",x"E5",x"CD",x"C9",x"0B",x"F1",x"33", -- 0x0D50
		x"21",x"54",x"13",x"E5",x"21",x"60",x"5D",x"E5", -- 0x0D58
		x"CD",x"7C",x"08",x"F1",x"F1",x"7D",x"B7",x"20", -- 0x0D60
		x"0D",x"3E",x"02",x"F5",x"33",x"21",x"60",x"13", -- 0x0D68
		x"E5",x"CD",x"C9",x"0B",x"F1",x"33",x"21",x"6C", -- 0x0D70
		x"5D",x"E5",x"21",x"60",x"5D",x"E5",x"CD",x"C7", -- 0x0D78
		x"0A",x"F1",x"F1",x"7D",x"B7",x"20",x"0D",x"3E", -- 0x0D80
		x"04",x"F5",x"33",x"21",x"95",x"13",x"E5",x"CD", -- 0x0D88
		x"C9",x"0B",x"F1",x"33",x"2A",x"74",x"5D",x"22", -- 0x0D90
		x"6D",x"5F",x"2A",x"76",x"5D",x"22",x"6F",x"5F", -- 0x0D98
		x"ED",x"4B",x"6D",x"5F",x"2A",x"6D",x"5F",x"11", -- 0x0DA0
		x"FF",x"FF",x"19",x"22",x"6D",x"5F",x"78",x"B1", -- 0x0DA8
		x"28",x"20",x"21",x"6C",x"5D",x"E5",x"21",x"60", -- 0x0DB0
		x"5D",x"E5",x"CD",x"C7",x"0A",x"F1",x"F1",x"7D", -- 0x0DB8
		x"B7",x"20",x"DD",x"3E",x"04",x"F5",x"33",x"21", -- 0x0DC0
		x"95",x"13",x"E5",x"CD",x"C9",x"0B",x"F1",x"33", -- 0x0DC8
		x"18",x"CE",x"11",x"00",x"60",x"ED",x"4B",x"6F", -- 0x0DD0
		x"5F",x"21",x"6F",x"5F",x"7E",x"C6",x"FF",x"77", -- 0x0DD8
		x"23",x"7E",x"CE",x"FF",x"77",x"78",x"B1",x"28", -- 0x0DE0
		x"25",x"D5",x"D5",x"21",x"60",x"5D",x"E5",x"CD", -- 0x0DE8
		x"C7",x"0A",x"F1",x"F1",x"7D",x"D1",x"B7",x"20", -- 0x0DF0
		x"0F",x"D5",x"3E",x"05",x"F5",x"33",x"21",x"AD", -- 0x0DF8
		x"13",x"E5",x"CD",x"C9",x"0B",x"F1",x"33",x"D1", -- 0x0E00
		x"ED",x"35",x"00",x"02",x"18",x"C7",x"3E",x"FF", -- 0x0E08
		x"D3",x"E7",x"C3",x"00",x"60",x"3E",x"FF",x"D3", -- 0x0E10
		x"E7",x"ED",x"91",x"10",x"81",x"21",x"64",x"00", -- 0x0E18
		x"CD",x"2E",x"03",x"3E",x"06",x"F5",x"33",x"21", -- 0x0E20
		x"C9",x"13",x"E5",x"CD",x"C9",x"0B",x"F1",x"33", -- 0x0E28
		x"C9",x"ED",x"91",x"43",x"00",x"ED",x"91",x"40", -- 0x0E30
		x"00",x"0E",x"00",x"79",x"D6",x"10",x"28",x"0E", -- 0x0E38
		x"06",x"00",x"21",x"E6",x"13",x"09",x"6E",x"7D", -- 0x0E40
		x"ED",x"92",x"41",x"0C",x"18",x"ED",x"0E",x"00", -- 0x0E48
		x"79",x"D6",x"10",x"C8",x"06",x"00",x"21",x"F6", -- 0x0E50
		x"13",x"09",x"6E",x"7D",x"ED",x"92",x"41",x"0C", -- 0x0E58
		x"18",x"EE",x"DD",x"E5",x"DD",x"21",x"00",x"00", -- 0x0E60
		x"DD",x"39",x"DD",x"7E",x"04",x"E6",x"1F",x"32", -- 0x0E68
		x"71",x"5F",x"DD",x"7E",x"05",x"21",x"72",x"5F", -- 0x0E70
		x"77",x"3E",x"17",x"96",x"30",x"02",x"36",x"17", -- 0x0E78
		x"DD",x"E1",x"C9",x"DD",x"E5",x"DD",x"21",x"00", -- 0x0E80
		x"00",x"DD",x"39",x"01",x"2B",x"10",x"DD",x"7E", -- 0x0E88
		x"04",x"1E",x"00",x"C6",x"E0",x"6F",x"7B",x"CE", -- 0x0E90
		x"FF",x"67",x"29",x"29",x"29",x"09",x"EB",x"2A", -- 0x0E98
		x"71",x"5F",x"3A",x"71",x"5F",x"6F",x"E5",x"CD", -- 0x0EA0
		x"8B",x"00",x"0E",x"00",x"79",x"D6",x"08",x"28", -- 0x0EA8
		x"0A",x"1A",x"13",x"77",x"ED",x"34",x"00",x"01", -- 0x0EB0
		x"0C",x"18",x"F1",x"21",x"71",x"5F",x"34",x"DD", -- 0x0EB8
		x"E1",x"C9",x"DD",x"E5",x"DD",x"21",x"00",x"00", -- 0x0EC0
		x"DD",x"39",x"DD",x"4E",x"04",x"DD",x"46",x"05", -- 0x0EC8
		x"0A",x"B7",x"28",x"0B",x"03",x"C5",x"F5",x"33", -- 0x0ED0
		x"CD",x"83",x"0E",x"33",x"C1",x"18",x"F1",x"DD", -- 0x0ED8
		x"E1",x"C9",x"3E",x"FF",x"D3",x"E7",x"06",x"0A", -- 0x0EE0
		x"3E",x"FF",x"D3",x"EB",x"10",x"FA",x"3E",x"FE", -- 0x0EE8
		x"D3",x"E7",x"3E",x"4C",x"CD",x"E7",x"0F",x"06", -- 0x0EF0
		x"09",x"DB",x"EB",x"10",x"FC",x"06",x"10",x"3E", -- 0x0EF8
		x"40",x"11",x"00",x"00",x"C5",x"CD",x"C1",x"0F", -- 0x0F00
		x"C1",x"D2",x"15",x"0F",x"10",x"F1",x"2E",x"00", -- 0x0F08
		x"3E",x"FF",x"D3",x"E7",x"C9",x"3E",x"48",x"11", -- 0x0F10
		x"AA",x"01",x"CD",x"CE",x"0F",x"21",x"A5",x"0F", -- 0x0F18
		x"38",x"03",x"21",x"B3",x"0F",x"01",x"78",x"00", -- 0x0F20
		x"C5",x"CD",x"3C",x"0F",x"C1",x"D2",x"3D",x"0F", -- 0x0F28
		x"10",x"F6",x"0D",x"20",x"F3",x"2E",x"00",x"3E", -- 0x0F30
		x"FF",x"D3",x"E7",x"C9",x"E9",x"3E",x"7A",x"11", -- 0x0F38
		x"00",x"00",x"CD",x"CE",x"0F",x"DA",x"35",x"0F", -- 0x0F40
		x"78",x"E6",x"40",x"32",x"73",x"5F",x"CC",x"60", -- 0x0F48
		x"0F",x"3E",x"FF",x"D3",x"E7",x"3A",x"73",x"5F", -- 0x0F50
		x"2E",x"03",x"FE",x"40",x"C8",x"2E",x"02",x"C9", -- 0x0F58
		x"3E",x"50",x"01",x"00",x"00",x"11",x"00",x"02", -- 0x0F60
		x"C3",x"AC",x"0F",x"E1",x"D1",x"C1",x"E3",x"3E", -- 0x0F68
		x"FE",x"D3",x"E7",x"3A",x"73",x"5F",x"B7",x"CC", -- 0x0F70
		x"99",x"0F",x"3E",x"51",x"CD",x"AC",x"0F",x"30", -- 0x0F78
		x"03",x"2E",x"00",x"C9",x"CD",x"0E",x"10",x"38", -- 0x0F80
		x"F8",x"01",x"EB",x"00",x"ED",x"B2",x"ED",x"B2", -- 0x0F88
		x"00",x"DB",x"EB",x"00",x"DB",x"EB",x"2E",x"01", -- 0x0F90
		x"C9",x"41",x"4A",x"53",x"1E",x"00",x"CB",x"22", -- 0x0F98
		x"CB",x"11",x"CB",x"10",x"C9",x"3E",x"41",x"01", -- 0x0FA0
		x"00",x"00",x"50",x"59",x"CD",x"E7",x"0F",x"B7", -- 0x0FA8
		x"C8",x"37",x"C9",x"3E",x"77",x"CD",x"A7",x"0F", -- 0x0FB0
		x"3E",x"69",x"01",x"00",x"40",x"51",x"59",x"18", -- 0x0FB8
		x"EB",x"01",x"00",x"00",x"CD",x"E7",x"0F",x"47", -- 0x0FC0
		x"E6",x"FE",x"78",x"20",x"E4",x"C9",x"CD",x"C1", -- 0x0FC8
		x"0F",x"D8",x"F5",x"CD",x"1C",x"10",x"67",x"CD", -- 0x0FD0
		x"1C",x"10",x"6F",x"CD",x"1C",x"10",x"57",x"CD", -- 0x0FD8
		x"1C",x"10",x"5F",x"44",x"4D",x"F1",x"C9",x"D3", -- 0x0FE0
		x"EB",x"F5",x"78",x"00",x"D3",x"EB",x"79",x"00", -- 0x0FE8
		x"D3",x"EB",x"7A",x"00",x"D3",x"EB",x"7B",x"00", -- 0x0FF0
		x"D3",x"EB",x"F1",x"FE",x"40",x"06",x"95",x"28", -- 0x0FF8
		x"08",x"FE",x"48",x"06",x"87",x"28",x"02",x"06", -- 0x1000
		x"FF",x"78",x"D3",x"EB",x"18",x"0E",x"06",x"0A", -- 0x1008
		x"C5",x"CD",x"1C",x"10",x"C1",x"FE",x"FE",x"C8", -- 0x1010
		x"10",x"F6",x"37",x"C9",x"01",x"64",x"00",x"DB", -- 0x1018
		x"EB",x"FE",x"FF",x"C0",x"10",x"F9",x"0D",x"20", -- 0x1020
		x"F6",x"C9",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1028
		x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10", -- 0x1030
		x"00",x"10",x"00",x"00",x"24",x"24",x"00",x"00", -- 0x1038
		x"00",x"00",x"00",x"00",x"24",x"7E",x"24",x"24", -- 0x1040
		x"7E",x"24",x"00",x"00",x"08",x"3E",x"28",x"3E", -- 0x1048
		x"0A",x"3E",x"08",x"00",x"62",x"64",x"08",x"10", -- 0x1050
		x"26",x"46",x"00",x"00",x"10",x"28",x"10",x"2A", -- 0x1058
		x"44",x"3A",x"00",x"00",x"08",x"10",x"00",x"00", -- 0x1060
		x"00",x"00",x"00",x"00",x"04",x"08",x"08",x"08", -- 0x1068
		x"08",x"04",x"00",x"00",x"20",x"10",x"10",x"10", -- 0x1070
		x"10",x"20",x"00",x"00",x"00",x"14",x"08",x"3E", -- 0x1078
		x"08",x"14",x"00",x"00",x"00",x"08",x"08",x"3E", -- 0x1080
		x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1088
		x"08",x"08",x"10",x"00",x"00",x"00",x"00",x"3E", -- 0x1090
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1098
		x"18",x"18",x"00",x"00",x"00",x"02",x"04",x"08", -- 0x10A0
		x"10",x"20",x"00",x"00",x"3C",x"46",x"4A",x"52", -- 0x10A8
		x"62",x"3C",x"00",x"00",x"18",x"28",x"08",x"08", -- 0x10B0
		x"08",x"3E",x"00",x"00",x"3C",x"42",x"02",x"3C", -- 0x10B8
		x"40",x"7E",x"00",x"00",x"3C",x"42",x"0C",x"02", -- 0x10C0
		x"42",x"3C",x"00",x"00",x"08",x"18",x"28",x"48", -- 0x10C8
		x"7E",x"08",x"00",x"00",x"7E",x"40",x"7C",x"02", -- 0x10D0
		x"42",x"3C",x"00",x"00",x"3C",x"40",x"7C",x"42", -- 0x10D8
		x"42",x"3C",x"00",x"00",x"7E",x"02",x"04",x"08", -- 0x10E0
		x"10",x"10",x"00",x"00",x"3C",x"42",x"3C",x"42", -- 0x10E8
		x"42",x"3C",x"00",x"00",x"3C",x"42",x"42",x"3E", -- 0x10F0
		x"02",x"3C",x"00",x"00",x"00",x"00",x"10",x"00", -- 0x10F8
		x"00",x"10",x"00",x"00",x"00",x"10",x"00",x"00", -- 0x1100
		x"10",x"10",x"20",x"00",x"00",x"04",x"08",x"10", -- 0x1108
		x"08",x"04",x"00",x"00",x"00",x"00",x"3E",x"00", -- 0x1110
		x"3E",x"00",x"00",x"00",x"00",x"10",x"08",x"04", -- 0x1118
		x"08",x"10",x"00",x"00",x"3C",x"42",x"04",x"08", -- 0x1120
		x"00",x"08",x"00",x"00",x"3C",x"4A",x"56",x"5E", -- 0x1128
		x"40",x"3C",x"00",x"00",x"3C",x"42",x"42",x"7E", -- 0x1130
		x"42",x"42",x"00",x"00",x"7C",x"42",x"7C",x"42", -- 0x1138
		x"42",x"7C",x"00",x"00",x"3C",x"42",x"40",x"40", -- 0x1140
		x"42",x"3C",x"00",x"00",x"78",x"44",x"42",x"42", -- 0x1148
		x"44",x"78",x"00",x"00",x"7E",x"40",x"7C",x"40", -- 0x1150
		x"40",x"7E",x"00",x"00",x"7E",x"40",x"7C",x"40", -- 0x1158
		x"40",x"40",x"00",x"00",x"3C",x"42",x"40",x"4E", -- 0x1160
		x"42",x"3C",x"00",x"00",x"42",x"42",x"7E",x"42", -- 0x1168
		x"42",x"42",x"00",x"00",x"3E",x"08",x"08",x"08", -- 0x1170
		x"08",x"3E",x"00",x"00",x"02",x"02",x"02",x"42", -- 0x1178
		x"42",x"3C",x"00",x"00",x"44",x"48",x"70",x"48", -- 0x1180
		x"44",x"42",x"00",x"00",x"40",x"40",x"40",x"40", -- 0x1188
		x"40",x"7E",x"00",x"00",x"42",x"66",x"5A",x"42", -- 0x1190
		x"42",x"42",x"00",x"00",x"42",x"62",x"52",x"4A", -- 0x1198
		x"46",x"42",x"00",x"00",x"3C",x"42",x"42",x"42", -- 0x11A0
		x"42",x"3C",x"00",x"00",x"7C",x"42",x"42",x"7C", -- 0x11A8
		x"40",x"40",x"00",x"00",x"3C",x"42",x"42",x"52", -- 0x11B0
		x"4A",x"3C",x"00",x"00",x"7C",x"42",x"42",x"7C", -- 0x11B8
		x"44",x"42",x"00",x"00",x"3C",x"40",x"3C",x"02", -- 0x11C0
		x"42",x"3C",x"00",x"00",x"FE",x"10",x"10",x"10", -- 0x11C8
		x"10",x"10",x"00",x"00",x"42",x"42",x"42",x"42", -- 0x11D0
		x"42",x"3C",x"00",x"00",x"42",x"42",x"42",x"42", -- 0x11D8
		x"24",x"18",x"00",x"00",x"42",x"42",x"42",x"42", -- 0x11E0
		x"5A",x"24",x"00",x"00",x"42",x"24",x"18",x"18", -- 0x11E8
		x"24",x"42",x"00",x"00",x"82",x"44",x"28",x"10", -- 0x11F0
		x"10",x"10",x"00",x"00",x"7E",x"04",x"08",x"10", -- 0x11F8
		x"20",x"7E",x"00",x"00",x"0E",x"08",x"08",x"08", -- 0x1200
		x"08",x"0E",x"00",x"00",x"00",x"40",x"20",x"10", -- 0x1208
		x"08",x"04",x"00",x"00",x"70",x"10",x"10",x"10", -- 0x1210
		x"10",x"70",x"00",x"00",x"10",x"38",x"54",x"10", -- 0x1218
		x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1220
		x"00",x"00",x"FF",x"00",x"1C",x"22",x"78",x"20", -- 0x1228
		x"20",x"7E",x"00",x"00",x"00",x"38",x"04",x"3C", -- 0x1230
		x"44",x"3C",x"00",x"00",x"20",x"20",x"3C",x"22", -- 0x1238
		x"22",x"3C",x"00",x"00",x"00",x"1C",x"20",x"20", -- 0x1240
		x"20",x"1C",x"00",x"00",x"04",x"04",x"3C",x"44", -- 0x1248
		x"44",x"3C",x"00",x"00",x"00",x"38",x"44",x"78", -- 0x1250
		x"40",x"3C",x"00",x"00",x"0C",x"10",x"18",x"10", -- 0x1258
		x"10",x"10",x"00",x"00",x"00",x"3C",x"44",x"44", -- 0x1260
		x"3C",x"04",x"38",x"00",x"40",x"40",x"78",x"44", -- 0x1268
		x"44",x"44",x"00",x"00",x"10",x"00",x"30",x"10", -- 0x1270
		x"10",x"38",x"00",x"00",x"04",x"00",x"04",x"04", -- 0x1278
		x"04",x"24",x"18",x"00",x"20",x"28",x"30",x"30", -- 0x1280
		x"28",x"24",x"00",x"00",x"10",x"10",x"10",x"10", -- 0x1288
		x"10",x"0C",x"00",x"00",x"00",x"68",x"54",x"54", -- 0x1290
		x"54",x"54",x"00",x"00",x"00",x"78",x"44",x"44", -- 0x1298
		x"44",x"44",x"00",x"00",x"00",x"38",x"44",x"44", -- 0x12A0
		x"44",x"38",x"00",x"00",x"00",x"78",x"44",x"44", -- 0x12A8
		x"78",x"40",x"40",x"00",x"00",x"3C",x"44",x"44", -- 0x12B0
		x"3C",x"04",x"06",x"00",x"00",x"1C",x"20",x"20", -- 0x12B8
		x"20",x"20",x"00",x"00",x"00",x"38",x"40",x"38", -- 0x12C0
		x"04",x"78",x"00",x"00",x"10",x"38",x"10",x"10", -- 0x12C8
		x"10",x"0C",x"00",x"00",x"00",x"44",x"44",x"44", -- 0x12D0
		x"44",x"38",x"00",x"00",x"00",x"44",x"44",x"28", -- 0x12D8
		x"28",x"10",x"00",x"00",x"00",x"44",x"54",x"54", -- 0x12E0
		x"54",x"28",x"00",x"00",x"00",x"44",x"28",x"10", -- 0x12E8
		x"28",x"44",x"00",x"00",x"00",x"44",x"44",x"44", -- 0x12F0
		x"3C",x"04",x"38",x"00",x"00",x"7C",x"08",x"10", -- 0x12F8
		x"20",x"7C",x"00",x"00",x"0E",x"08",x"30",x"08", -- 0x1300
		x"08",x"0E",x"00",x"00",x"08",x"08",x"08",x"08", -- 0x1308
		x"08",x"08",x"00",x"00",x"70",x"10",x"0C",x"10", -- 0x1310
		x"10",x"70",x"00",x"00",x"14",x"28",x"00",x"00", -- 0x1318
		x"00",x"00",x"00",x"3C",x"42",x"99",x"A1",x"A1", -- 0x1320
		x"99",x"42",x"3C",x"46",x"41",x"54",x"31",x"36", -- 0x1328
		x"20",x"20",x"20",x"00",x"46",x"41",x"54",x"33", -- 0x1330
		x"32",x"20",x"20",x"20",x"00",x"45",x"72",x"72", -- 0x1338
		x"6F",x"72",x"20",x"4D",x"6F",x"75",x"6E",x"74", -- 0x1340
		x"69",x"6E",x"67",x"20",x"53",x"44",x"20",x"43", -- 0x1348
		x"61",x"72",x"64",x"00",x"54",x"42",x"42",x"4C", -- 0x1350
		x"55",x"45",x"20",x"20",x"46",x"57",x"20",x"00", -- 0x1358
		x"54",x"42",x"42",x"4C",x"55",x"45",x"2E",x"46", -- 0x1360
		x"57",x"20",x"4E",x"6F",x"74",x"20",x"46",x"6F", -- 0x1368
		x"75",x"6E",x"64",x"00",x"54",x"42",x"42",x"4C", -- 0x1370
		x"55",x"45",x"20",x"20",x"54",x"42",x"55",x"00", -- 0x1378
		x"54",x"42",x"42",x"4C",x"55",x"45",x"2E",x"54", -- 0x1380
		x"42",x"55",x"20",x"4E",x"6F",x"74",x"20",x"46", -- 0x1388
		x"6F",x"75",x"6E",x"64",x"00",x"45",x"72",x"72", -- 0x1390
		x"6F",x"72",x"20",x"52",x"65",x"61",x"64",x"69", -- 0x1398
		x"6E",x"67",x"20",x"54",x"42",x"42",x"4C",x"55", -- 0x13A0
		x"45",x"2E",x"46",x"57",x"00",x"45",x"72",x"72", -- 0x13A8
		x"6F",x"72",x"20",x"4C",x"6F",x"61",x"64",x"69", -- 0x13B0
		x"6E",x"67",x"20",x"55",x"50",x"44",x"41",x"54", -- 0x13B8
		x"45",x"20",x"4D",x"6F",x"64",x"75",x"6C",x"65", -- 0x13C0
		x"00",x"46",x"61",x"69",x"6C",x"65",x"64",x"20", -- 0x13C8
		x"74",x"6F",x"20",x"53",x"74",x"61",x"72",x"74", -- 0x13D0
		x"20",x"5A",x"58",x"20",x"4E",x"65",x"78",x"74", -- 0x13D8
		x"20",x"43",x"6F",x"72",x"65",x"00",x"00",x"02", -- 0x13E0
		x"A0",x"A2",x"14",x"16",x"B4",x"B6",x"00",x"03", -- 0x13E8
		x"E0",x"E7",x"1C",x"1F",x"FC",x"FF",x"00",x"02", -- 0x13F0
		x"A0",x"A2",x"14",x"16",x"B4",x"B6",x"00",x"03", -- 0x13F8
		x"E0",x"E7",x"1C",x"1F",x"FC",x"FF",x"FF",x"FF", -- 0x1400
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1408
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1410
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1418
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1420
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1428
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1430
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1438
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1440
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1448
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1450
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1458
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1460
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1468
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1470
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1480
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1488
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1490
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1498
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1500
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1508
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1510
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1520
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1528
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1530
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1538
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1540
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1548
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1550
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1558
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1560
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1568
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1570
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1578
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1580
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1588
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1590
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1598
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1600
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1608
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1610
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1618
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1620
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1628
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1630
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1640
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1658
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1660
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1668
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1680
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1688
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1690
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1698
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1700
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1708
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1710
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1718
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1720
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1728
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1730
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1738
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1740
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1748
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1750
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1758
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1760
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1768
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1788
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1790
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1800
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1808
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1810
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1818
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1820
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1828
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1830
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1838
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1840
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1848
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1850
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1858
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1860
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1868
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1870
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1878
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1880
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1888
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1890
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1898
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1900
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1908
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1910
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1918
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1920
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1928
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1930
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1938
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1940
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1948
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1950
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1958
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1960
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1968
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1978
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1980
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1988
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1990
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1998
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1ED8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x1FF8
	);

begin

	process(clk)
	begin
		if rising_edge(clk) then
			data <= ROM(to_integer(unsigned(addr)));
		end if;
	end process;
end RTL;
